module counter (  input clk,
                  input rstn,
                  output reg[3:0] out);
endmodule

module counter2 (  input clk,
                  input rstn,
                  output reg[3:0] out);
endmodule